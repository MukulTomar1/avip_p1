`ifndef GLOBALS_PKG_INCLUDED_
`define GLOBALS_PKG_INCLUDED_

//--------------------------------------------------------------------------------------------
// global pkg for all variables 
//--------------------------------------------------------------------------------------------

package globals_pkg;

// NO_OF_SLAVES to be connected to the spi_interface

parameter int NO_OF_SLAVES = 1;

endpackage : globals_pkg 

`endif

