module hvl_top;

  import test_pkg::*;
  import uvm_pkg::*;


  initial
  begin
    run_test("base_test");
  end

endmodule : hvl_top
