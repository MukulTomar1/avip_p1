`ifndef P_IF_INCLUDED_
`define P_IF_INCLUDED_
//--------------------------------------------------------------------------------------------
// Module       : Interface
// Description  : Declaration of pin level signals as logic
//--------------------------------------------------------------------------------------------
interface p_if;

//--------------------------------------------------------------------------------------------
// mention all the signals here
//--------------------------------------------------------------------------------------------


endinterface : p_if

`endif
